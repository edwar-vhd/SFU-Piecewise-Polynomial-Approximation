library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity LUT_C1_ln2 is
	generic(
		word_bits	:natural:=19;
		bus_bits	:natural:=20;
		add_bits	:natural:=7
	);
	port(
		addr		:in std_logic_vector(add_bits-1 downto 0);
		data		:out std_logic_vector(bus_bits-1 downto 0)
	);
end entity;

architecture behav of LUT_C1_ln2 is
	type storage is array (0 to 2**add_bits-1) of std_logic_vector(word_bits-1 downto 0);
	signal rom:storage:=(
		"1011100010101001000",
		"1011011100111011000",
		"1011010111010010000",
		"1011010001101111000",
		"1011001100010001000",
		"1011000110111000000",
		"1011000001100101000",
		"1010111100010110000",
		"1010110111001100000",
		"1010110010001000000",
		"1010101101001000000",
		"1010101000001100000",
		"1010100011010101000",
		"1010011110100011000",
		"1010011001110100000",
		"1010010101001011000",
		"1010010000100101000",
		"1010001100000011000",
		"1010000111100101000",
		"1010000011001011000",
		"1001111110110101000",
		"1001111010100011000",
		"1001110110010100000",
		"1001110010001001000",
		"1001101110000001000",
		"1001101001111101000",
		"1001100101111100000",
		"1001100001111111000",
		"1001011110000100000",
		"1001011010001101000",
		"1001010110011001000",
		"1001010010101000000",
		"1001001110111011000",
		"1001001011010000000",
		"1001000111101000000",
		"1001000100000011000",
		"1001000000100000000",
		"1000111101000001000",
		"1000111001100100000",
		"1000110110001001000",
		"1000110010110010000",
		"1000101111011101000",
		"1000101100001010000",
		"1000101000111010000",
		"1000100101101100000",
		"1000100010100001000",
		"1000011111011000000",
		"1000011100010001000",
		"1000011001001101000",
		"1000010110001010000",
		"1000010011001010000",
		"1000010000001100000",
		"1000001101010001000",
		"1000001010010111000",
		"1000000111011111000",
		"1000000100101001000",
		"1000000001110110000",
		"0111111111000100000",
		"0111111100010100000",
		"0111111001100110000",
		"0111110110111010000",
		"0111110100010000000",
		"0111110001100111000",
		"0111101111000000000",
		"0111101100011011000",
		"0111101001111000000",
		"0111100111010111000",
		"0111100100110111000",
		"0111100010011000000",
		"0111011111111100000",
		"0111011101100000000",
		"0111011011000111000",
		"0111011000101111000",
		"0111010110011000000",
		"0111010100000011000",
		"0111010001110000000",
		"0111001111011110000",
		"0111001101001101000",
		"0111001010111110000",
		"0111001000110000000",
		"0111000110100011000",
		"0111000100011000000",
		"0111000010001110000",
		"0111000000000110000",
		"0110111101111110000",
		"0110111011111000000",
		"0110111001110100000",
		"0110110111110000000",
		"0110110101101110000",
		"0110110011101101000",
		"0110110001101101000",
		"0110101111101110000",
		"0110101101110000000",
		"0110101011110100000",
		"0110101001111001000",
		"0110100111111110000",
		"0110100110000101000",
		"0110100100001101000",
		"0110100010010110000",
		"0110100000100000000",
		"0110011110101011000",
		"0110011100110111000",
		"0110011011000101000",
		"0110011001010011000",
		"0110010111100010000",
		"0110010101110010000",
		"0110010100000011000",
		"0110010010010101000",
		"0110010000101000000",
		"0110001110111011000",
		"0110001101010000000",
		"0110001011100110000",
		"0110001001111100000",
		"0110001000010100000",
		"0110000110101100000",
		"0110000101000101000",
		"0110000011011111000",
		"0110000001111010000",
		"0110000000010101000",
		"0101111110110010000",
		"0101111101001111000",
		"0101111011101101000",
		"0101111010001100000",
		"0101111000101011000",
		"0101110111001100000",
		"0101110101101101000",
		"0101110100001111000",
		"0101110010110001000"
	);
begin
	data <= "0"&rom(to_integer(unsigned(addr)));
end architecture;