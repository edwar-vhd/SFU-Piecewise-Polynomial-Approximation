library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity LUT_C0_exp is
	generic(
		word_bits	:natural:=25;
		bus_bits	:natural:=29;
		add_bits	:natural:=6
	);
	port(
		addr		:in std_logic_vector(add_bits-1 downto 0);
		data		:out std_logic_vector(bus_bits-1 downto 0)
	);
end entity;

architecture behav of LUT_C0_exp is
	type storage is array (0 to 2**add_bits-1) of std_logic_vector(word_bits-1 downto 0);
	signal rom:storage:=(
		"0000000000000000000000000",
		"0000001011001001101001000",
		"0000010110011011000011010",
		"0000100001110100010100011",
		"0000101101010101100001101",
		"0000111000111110110000110",
		"0001000100110000000111010",
		"0001010000101001101010110",
		"0001011100101011100000111",
		"0001101000110101101111101",
		"0001110101001000011100110",
		"0010000001100011101110001",
		"0010001110000111101001110",
		"0010011010110100010101101",
		"0010100111101001110111110",
		"0010110100101000010110101",
		"0011000001101111111000001",
		"0011001111000000100010110",
		"0011011100011010011100111",
		"0011101001111101101100110",
		"0011110111101010011001001",
		"0100000101100000101000100",
		"0100010011100000100001100",
		"0100100001101010001010111",
		"0100101111111101101011010",
		"0100111110011011001001111",
		"0101001101000010101101011",
		"0101011011110100011100111",
		"0101101010110000011111011",
		"0101111001110110111100011",
		"0110001001000111111010110",
		"0110011000100011100010000",
		"0110101000001001111001101",
		"0110110111111011001000111",
		"0111000111110111010111101",
		"0111010111111110101101011",
		"0111101000010001010001110",
		"0111111000101111001100111",
		"1000001001011000100110011",
		"1000011010001101100110011",
		"1000101011001110010101000",
		"1000111100011010111010011",
		"1001001101110011011110110",
		"1001011111011000001010100",
		"1001110001001001000110000",
		"1010000011000110011001111",
		"1010010101010000001110110",
		"1010100111100110101101011",
		"1010111010001001111110011",
		"1011001100111010001010111",
		"1011011111110111011011110",
		"1011110011000001111010010",
		"1100000110011001101111100",
		"1100011001111111000100110",
		"1100101101110010000011100",
		"1101000001110010110101001",
		"1101010110000001100011100",
		"1101101010011110011000000",
		"1101111111001001011100110",
		"1110010100000010111011101",
		"1110101001001010111110100",
		"1110111110100001101111110",
		"1111010100000111011001011",
		"1111101001111100000110000"
	);
begin
	data <= "01"&rom(to_integer(unsigned(addr)))&"00";
end architecture;