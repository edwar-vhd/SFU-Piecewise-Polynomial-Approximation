library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity LUT_C0_reci_sqrt_2_4 is
	generic(
		word_bits	:natural:=24;
		bus_bits	:natural:=29;
		add_bits	:natural:=7
	);
	port(
		addr		:in std_logic_vector(add_bits-1 downto 0);
		data		:out std_logic_vector(bus_bits-1 downto 0)
	);
end entity;

architecture behav of LUT_C0_reci_sqrt_2_4 is
	type storage is array (0 to 2**add_bits-1) of std_logic_vector(word_bits-1 downto 0);
	signal rom:storage:=(
		"110101000001001111001100",
		"110100010100001111101111",
		"110011100111110001100101",
		"110010111011110100000101",
		"110010010000010110100110",
		"110001100101011000100011",
		"110000111010111001010110",
		"110000010000111000011010",
		"101111100111010101001100",
		"101110111110001111001001",
		"101110010101100101101110",
		"101101101101011000011100",
		"101101000101100110110001",
		"101100011110010000001110",
		"101011110111010100010101",
		"101011010000110010101000",
		"101010101010101010101010",
		"101010000100111011111110",
		"101001011111100110001000",
		"101000111010101000101110",
		"101000010110000011010100",
		"100111110001110101100010",
		"100111001101111110111110",
		"100110101010011111001111",
		"100110000111010101111101",
		"100101100100100010110000",
		"100101000010000101010010",
		"100100011111111101001101",
		"100011111110001010001001",
		"100011011100101011110011",
		"100010111011100001110100",
		"100010011010101011111000",
		"100001111010001001101100",
		"100001011001111010111011",
		"100000111001111111010010",
		"100000011010010110011111",
		"011111111011000000001110",
		"011111011011111100001111",
		"011110111101001010001111",
		"011110011110101001111110",
		"011110000000011011001010",
		"011101100010011101100010",
		"011101000100110000110111",
		"011100100111010100111000",
		"011100001010001001010111",
		"011011101101001110000011",
		"011011010000100010101110",
		"011010110100000111001010",
		"011010010111111011000111",
		"011001111011111110011000",
		"011001100000010000110000",
		"011001000100110001111111",
		"011000101001100001111011",
		"011000001110100000010100",
		"010111110011101100111111",
		"010111011001000111101111",
		"010110111110110000011000",
		"010110100100100110101110",
		"010110001010101010100101",
		"010101110000111011110001",
		"010101010111011010000111",
		"010100111110000101011100",
		"010100100100111101100101",
		"010100001100000010010111",
		"010011110011010011101000",
		"010011011010110001001101",
		"010011000010011010111101",
		"010010101010010000101100",
		"010010010010010010010010",
		"010001111010011111100100",
		"010001100010111000011010",
		"010001001011011100101001",
		"010000110100001100001010",
		"010000011101000110110010",
		"010000000110001100011001",
		"001111101111011100110110",
		"001111011000111000000010",
		"001111000010011101110010",
		"001110101100001110000000",
		"001110010110001000100011",
		"001110000000001101010011",
		"001101101010011100001001",
		"001101010100110100111100",
		"001100111111010111100101",
		"001100101010000011111101",
		"001100010100111001111100",
		"001011111111111001011011",
		"001011101011000010010100",
		"001011010110010100011110",
		"001011000001101111110100",
		"001010101101010100001110",
		"001010011001000001100110",
		"001010000100110111110101",
		"001001110000110110110101",
		"001001011100111110100000",
		"001001001001001110101111",
		"001000110101100111011100",
		"001000100010001000100010",
		"001000001110110001111001",
		"000111111011100011011101",
		"000111101000011101001000",
		"000111010101011110110100",
		"000111000010101000011011",
		"000110101111111001111000",
		"000110011101010011000110",
		"000110001010110011111110",
		"000101111000011100011101",
		"000101100110001100011100",
		"000101010100000011110111",
		"000101000010000010101001",
		"000100110000001000101100",
		"000100011110010101111100",
		"000100001100101010010100",
		"000011111011000101101111",
		"000011101001101000001001",
		"000011011000010001011101",
		"000011000111000001100110",
		"000010110101111000100000",
		"000010100100110110000111",
		"000010010011111010010110",
		"000010000011000101001000",
		"000001110010010110011011",
		"000001100001101110001001",
		"000001010001001100001111",
		"000001000000110000101000",
		"000000110000011011010001",
		"000000100000001100000101",
		"000000010000000011000000"
	);
begin
	data <= "0010"&rom(to_integer(unsigned(addr)))&"0";
end architecture;