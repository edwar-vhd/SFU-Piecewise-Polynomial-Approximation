library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity LUT_C0_sqrt_1_2 is
	generic(
		word_bits	:natural:=26;
		bus_bits	:natural:=29;
		add_bits	:natural:=6
	);
	port(
		addr		:in std_logic_vector(add_bits-1 downto 0);
		data		:out std_logic_vector(bus_bits-1 downto 0)
	);
end entity;

architecture behav of LUT_C0_sqrt_1_2 is
	type storage is array (0 to 2**add_bits-1) of std_logic_vector(word_bits-1 downto 0);
	signal rom:storage:=(
		"00000000000000000000000000",
		"00000011111111000000100000",
		"00000111111100000011111000",
		"00001011110111001101001000",
		"00001111110000011110110100",
		"00010011100111111011100100",
		"00010111011101100110000100",
		"00011011010001100000100100",
		"00011111000011101101100100",
		"00100010110100001111010100",
		"00100110100011000111111100",
		"00101010010000011001101000",
		"00101101111100000110011000",
		"00110001100110010000010000",
		"00110101001110111001001000",
		"00111000110110000010110100",
		"00111100011011101111001100",
		"01000000000000000000000000",
		"01000011100010110110111000",
		"01000111000100010101100000",
		"01001010100100011101011100",
		"01001110000011010000010000",
		"01010001100000101111011100",
		"01010100111100111100011100",
		"01011000010111111000101100",
		"01011011110001100101100000",
		"01011111001010000100010100",
		"01100010100001010110011000",
		"01100101110111011100111000",
		"01101001001100011001001100",
		"01101100100000001100011000",
		"01101111110010110111101000",
		"01110011000100011100001000",
		"01110110010100111010111100",
		"01111001100100010101001100",
		"01111100110010101011110100",
		"10000000000000000000000000",
		"10000011001100010010100100",
		"10000110010111100100101000",
		"10001001100001110111000000",
		"10001100101011001010101100",
		"10001111110011100000101000",
		"10010010111010111001101000",
		"10010110000001010110100100",
		"10011001000110111000010100",
		"10011100001011011111101100",
		"10011111001111001101011100",
		"10100010010010000010011000",
		"10100101010011111111010100",
		"10101000010101000100111100",
		"10101011010101010100000000",
		"10101110010100101101001100",
		"10110001010011010001010000",
		"10110100010001000000111000",
		"10110111001101111100101100",
		"10111010001010000101011000",
		"10111101000101011011101000",
		"11000000000000000000000000",
		"11000010111001110011000100",
		"11000101110010110101100100",
		"11001000101011001000000000",
		"11001011100010101011000000",
		"11001110011001011111000100",
		"11010001001111100100110100"
	);
begin
	data <= "010"&rom(to_integer(unsigned(addr)));
end architecture;