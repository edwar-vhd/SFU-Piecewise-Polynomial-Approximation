library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity LUT_C2_ln2e0 is
	generic(
		word_bits	:natural:=12;
		bus_bits	:natural:=14;
		add_bits	:natural:=6
	);
	port(
		addr		:in std_logic_vector(add_bits-1 downto 0);
		data		:out std_logic_vector(bus_bits-1 downto 0)
	);
end entity;

architecture behav of LUT_C2_ln2e0 is
	type storage is array (0 to 2**add_bits-1) of std_logic_vector(word_bits-1 downto 0);
	signal rom:storage:=(
		"111100011000",
		"111010011000",
		"111000011000",
		"110110100000",
		"110100110000",
		"110011000000",
		"110001011000",
		"101111111000",
		"101110011000",
		"101101000000",
		"101011101000",
		"101010011000",
		"101001001000",
		"100111111000",
		"100110110000",
		"100101101000",
		"100100101000",
		"100011100000",
		"100010101000",
		"100001101000",
		"100000110000",
		"011111111000",
		"011111000000",
		"011110010000",
		"011101100000",
		"011100110000",
		"011100000000",
		"011011010000",
		"011010101000",
		"011010000000",
		"011001011000",
		"011000110000",
		"011000001000",
		"010111101000",
		"010111000000",
		"010110100000",
		"010110000000",
		"010101100000",
		"010101000000",
		"010100100000",
		"010100001000",
		"010011101000",
		"010011010000",
		"010010110000",
		"010010011000",
		"010010000000",
		"010001101000",
		"010001010000",
		"010000111000",
		"010000101000",
		"010000010000",
		"001111111000",
		"001111101000",
		"001111010000",
		"001111000000",
		"001110110000",
		"001110011000",
		"001110001000",
		"001101111000",
		"001101101000",
		"001101011000",
		"001101001000",
		"001100111000",
		"001100101000"
	);
begin
	data <= "00"&rom(to_integer(unsigned(addr)));
end architecture;