library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity LUT_C2_sin is
	generic(
		word_bits	:natural:=12;
		bus_bits	:natural:=14;
		add_bits	:natural:=6
	);
	port(
		addr		:in std_logic_vector(add_bits-1 downto 0);
		data		:out std_logic_vector(bus_bits-1 downto 0)
	);
end entity;

architecture behav of LUT_C2_sin is
	type storage is array (0 to 2**add_bits-1) of std_logic_vector(word_bits-1 downto 0);
	signal rom:storage:=(
		"000000011111",
		"000001011111",
		"000010011111",
		"000011011111",
		"000100011111",
		"000101011111",
		"000110011111",
		"000111011110",
		"001000011110",
		"001001011101",
		"001010011100",
		"001011011100",
		"001100011010",
		"001101011001",
		"001110011000",
		"001111010110",
		"010000010100",
		"010001010010",
		"010010001111",
		"010011001100",
		"010100001001",
		"010101000110",
		"010110000010",
		"010110111110",
		"010111111001",
		"011000110101",
		"011001101111",
		"011010101010",
		"011011100100",
		"011100011101",
		"011101010110",
		"011110001111",
		"011111000111",
		"011111111111",
		"100000110110",
		"100001101101",
		"100010100011",
		"100011011000",
		"100100001110",
		"100101000010",
		"100101110110",
		"100110101001",
		"100111011100",
		"101000001110",
		"101000111111",
		"101001110000",
		"101010100000",
		"101011010000",
		"101011111111",
		"101100101101",
		"101101011010",
		"101110000111",
		"101110110011",
		"101111011110",
		"110000001001",
		"110000110011",
		"110001011100",
		"110010000100",
		"110010101011",
		"110011010010",
		"110011111000",
		"110100011101",
		"110101000001",
		"110101100101"
	);
begin
	data <= "10"&rom(to_integer(unsigned(addr)));
end architecture;