library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity LUT_C1_reci_sqrt_2_4 is
	generic(
		word_bits	:natural:=17;
		bus_bits	:natural:=20;
		add_bits	:natural:=7
	);
	port(
		addr		:in std_logic_vector(add_bits-1 downto 0);
		data		:out std_logic_vector(bus_bits-1 downto 0)
	);
end entity;

architecture behav of LUT_C1_reci_sqrt_2_4 is
	type storage is array (0 to 2**add_bits-1) of std_logic_vector(word_bits-1 downto 0);
	signal rom:storage:=(
		"10110101000000100",
		"10110010111010100",
		"10110000110110100",
		"10101110110101000",
		"10101100110110000",
		"10101010111001100",
		"10101000111111100",
		"10100111000111100",
		"10100101010001100",
		"10100011011110000",
		"10100001101100100",
		"10011111111101000",
		"10011110001111100",
		"10011100100100000",
		"10011010111010100",
		"10011001010010100",
		"10010111101100100",
		"10010110001000100",
		"10010100100110000",
		"10010011000101000",
		"10010001100101100",
		"10010000001000000",
		"10001110101100000",
		"10001101010001100",
		"10001011111000100",
		"10001010100000100",
		"10001001001010100",
		"10000111110101100",
		"10000110100010000",
		"10000101010000000",
		"10000011111111100",
		"10000010101111100",
		"10000001100001100",
		"10000000010100000",
		"01111111001000100",
		"01111101111101100",
		"01111100110100000",
		"01111011101011100",
		"01111010100100000",
		"01111001011101100",
		"01111000011000100",
		"01110111010100000",
		"01110110010001000",
		"01110101001110100",
		"01110100001101000",
		"01110011001101000",
		"01110010001101100",
		"01110001001110100",
		"01110000010001000",
		"01101111010100100",
		"01101110011000100",
		"01101101011101000",
		"01101100100011000",
		"01101011101001100",
		"01101010110000100",
		"01101001111001000",
		"01101001000001100",
		"01101000001011000",
		"01100111010101100",
		"01100110100000100",
		"01100101101100000",
		"01100100111000100",
		"01100100000101100",
		"01100011010011100",
		"01100010100010000",
		"01100001110001000",
		"01100001000000100",
		"01100000010001000",
		"01011111100010000",
		"01011110110011100",
		"01011110000101100",
		"01011101011000000",
		"01011100101011100",
		"01011011111111000",
		"01011011010011100",
		"01011010101000100",
		"01011001111101100",
		"01011001010011100",
		"01011000101010000",
		"01011000000001000",
		"01010111011000100",
		"01010110110000100",
		"01010110001000100",
		"01010101100001100",
		"01010100111011000",
		"01010100010100100",
		"01010011101111000",
		"01010011001001100",
		"01010010100100100",
		"01010010000000000",
		"01010001011100000",
		"01010000111000100",
		"01010000010101000",
		"01001111110010100",
		"01001111010000000",
		"01001110101110000",
		"01001110001100000",
		"01001101101010100",
		"01001101001010000",
		"01001100101001000",
		"01001100001001000",
		"01001011101001000",
		"01001011001001100",
		"01001010101010100",
		"01001010001011100",
		"01001001101101000",
		"01001001001110100",
		"01001000110001000",
		"01001000010011100",
		"01000111110110000",
		"01000111011001000",
		"01000110111100100",
		"01000110100000000",
		"01000110000100000",
		"01000101101000100",
		"01000101001101000",
		"01000100110001100",
		"01000100010110100",
		"01000011111100000",
		"01000011100001100",
		"01000011000111100",
		"01000010101101100",
		"01000010010100000",
		"01000001111010100",
		"01000001100001100",
		"01000001001001000",
		"01000000110000000",
		"01000000011000000"
	);
begin
	data <= "100"&rom(to_integer(unsigned(addr)));
end architecture;