library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity LUT_C0_exp is
	generic(
		word_bits	:natural:=27;
		bus_bits	:natural:=29;
		add_bits	:natural:=6
	);
	port(
		addr		:in std_logic_vector(add_bits-1 downto 0);
		data		:out std_logic_vector(bus_bits-1 downto 0)
	);
end entity;

architecture behav of LUT_C0_exp is
	type storage is array (0 to 2**add_bits-1) of std_logic_vector(word_bits-1 downto 0);
	signal rom:storage:=(
		"000000000000000000000000000",
		"000000101100100110100100000",
		"000001011001101100001101000",
		"000010000111010001010001100",
		"000010110101010110000110100",
		"000011100011111011000011000",
		"000100010011000000011101000",
		"000101000010100110101011000",
		"000101110010101110000011100",
		"000110100011010110111110100",
		"000111010100100001110011000",
		"001000000110001110111000100",
		"001000111000011110100111000",
		"001001101011010001010110100",
		"001010011110100111011111000",
		"001011010010100001011010100",
		"001100000110111111100000100",
		"001100111100000010001011000",
		"001101110001101001110011100",
		"001110100111110110110011000",
		"001111011110101001100100100",
		"010000010110000010100010000",
		"010001001110000010000110000",
		"010010000110101000101011100",
		"010010111111110110101101000",
		"010011111001101100100111100",
		"010100110100001010110101100",
		"010101101111010001110011100",
		"010110101011000001111101100",
		"010111100111011011110001100",
		"011000100100011111101011000",
		"011001100010001110001000000",
		"011010100000100111100110100",
		"011011011111101100100011100",
		"011100011111011101011110100",
		"011101011111111010110101100",
		"011110100001000101000111000",
		"011111100010111100110011100",
		"100000100101100010011001100",
		"100001101000110110011001100",
		"100010101100111001010100000",
		"100011110001101011101001100",
		"100100110111001101111011000",
		"100101111101100000101010000",
		"100111000100100100011000000",
		"101000001100011001100111100",
		"101001010101000000111011000",
		"101010011110011010110101100",
		"101011101000100111111001100",
		"101100110011101000101011100",
		"101101111111011101101111000",
		"101111001100000111101001000",
		"110000011001100110111110000",
		"110001100111111100010011000",
		"110010110111001000001110000",
		"110100000111001011010100100",
		"110101011000000110001110000",
		"110110101001111001100000000",
		"110111111100100101110011000",
		"111001010000001011101110100",
		"111010100100101011111010000",
		"111011111010000110111111000",
		"111101010000011101100101100",
		"111110100111110000011000000"
	);
begin
	data <= "01"&rom(to_integer(unsigned(addr)));
end architecture;