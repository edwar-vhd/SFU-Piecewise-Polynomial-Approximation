library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity LUT_C2_exp is
	generic(
		word_bits	:natural:=12;
		bus_bits	:natural:=14;
		add_bits	:natural:=6
	);
	port(
		addr		:in std_logic_vector(add_bits-1 downto 0);
		data		:out std_logic_vector(bus_bits-1 downto 0)
	);
end entity;

architecture behav of LUT_C2_exp is
	type storage is array (0 to 2**add_bits-1) of std_logic_vector(word_bits-1 downto 0);
	signal rom:storage:=(
		"011110111000",
		"011111010000",
		"011111100100",
		"011111111000",
		"100000010000",
		"100000101000",
		"100000111100",
		"100001010100",
		"100001101100",
		"100010000100",
		"100010011100",
		"100010110100",
		"100011001100",
		"100011100100",
		"100011111100",
		"100100010100",
		"100100110000",
		"100101001000",
		"100101100100",
		"100101111100",
		"100110011000",
		"100110110000",
		"100111001100",
		"100111101000",
		"101000000100",
		"101000100000",
		"101000111100",
		"101001011000",
		"101001110100",
		"101010010100",
		"101010110000",
		"101011010000",
		"101011101100",
		"101100001100",
		"101100101000",
		"101101001000",
		"101101101000",
		"101110001000",
		"101110101000",
		"101111001000",
		"101111101000",
		"110000001100",
		"110000101100",
		"110001010000",
		"110001110000",
		"110010010100",
		"110010111000",
		"110011011000",
		"110011111100",
		"110100100000",
		"110101001000",
		"110101101100",
		"110110010000",
		"110110111000",
		"110111011100",
		"111000000100",
		"111000101100",
		"111001010100",
		"111001111100",
		"111010100100",
		"111011001100",
		"111011110100",
		"111100100000",
		"111101001000"
	);
begin
	data <= "00"&rom(to_integer(unsigned(addr)));
end architecture;