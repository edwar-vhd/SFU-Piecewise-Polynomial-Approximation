library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity LUT_C2_sqrt_1_2 is
	generic(
		word_bits	:natural:=10;
		bus_bits	:natural:=14;
		add_bits	:natural:=6
	);
	port(
		addr		:in std_logic_vector(add_bits-1 downto 0);
		data		:out std_logic_vector(bus_bits-1 downto 0)
	);
end entity;

architecture behav of LUT_C2_sqrt_1_2 is
	type storage is array (0 to 2**add_bits-1) of std_logic_vector(word_bits-1 downto 0);
	signal rom:storage:=(
		"1111110100",
		"1111011100",
		"1111000100",
		"1110110000",
		"1110011100",
		"1110001000",
		"1101110100",
		"1101100000",
		"1101010000",
		"1101000000",
		"1100101100",
		"1100011100",
		"1100001100",
		"1100000000",
		"1011110000",
		"1011100000",
		"1011010100",
		"1011001000",
		"1010111000",
		"1010101100",
		"1010100000",
		"1010010100",
		"1010001000",
		"1010000000",
		"1001110100",
		"1001101000",
		"1001100000",
		"1001010100",
		"1001001100",
		"1001000000",
		"1000111000",
		"1000110000",
		"1000101000",
		"1000100000",
		"1000011000",
		"1000010000",
		"1000001000",
		"1000000000",
		"0111111000",
		"0111110000",
		"0111101000",
		"0111100000",
		"0111011100",
		"0111010100",
		"0111001100",
		"0111001000",
		"0111000000",
		"0110111100",
		"0110110100",
		"0110110000",
		"0110101000",
		"0110100100",
		"0110100000",
		"0110011000",
		"0110010100",
		"0110010000",
		"0110001100",
		"0110000100",
		"0110000000",
		"0101111100",
		"0101111000",
		"0101110100",
		"0101110000",
		"0101101100"
	);
begin
	data <= "1000"&rom(to_integer(unsigned(addr)));
end architecture;