library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity LUT_C2_ln2 is
	generic(
		word_bits	:natural:=10;
		bus_bits	:natural:=14;
		add_bits	:natural:=7
	);
	port(
		addr		:in std_logic_vector(add_bits-1 downto 0);
		data		:out std_logic_vector(bus_bits-1 downto 0)
	);
end entity;

architecture behav of LUT_C2_ln2 is
	type storage is array (0 to 2**add_bits-1) of std_logic_vector(word_bits-1 downto 0);
	signal rom:storage:=(
		"1011011100",
		"1011010001",
		"1011000110",
		"1010111011",
		"1010110001",
		"1010100111",
		"1010011100",
		"1010010011",
		"1010001001",
		"1010000000",
		"1001110110",
		"1001101101",
		"1001100101",
		"1001011100",
		"1001010011",
		"1001001011",
		"1001000011",
		"1000111011",
		"1000110011",
		"1000101100",
		"1000100100",
		"1000011101",
		"1000010110",
		"1000001111",
		"1000001000",
		"1000000001",
		"0111111011",
		"0111110100",
		"0111101110",
		"0111100111",
		"0111100001",
		"0111011011",
		"0111010101",
		"0111010000",
		"0111001010",
		"0111000100",
		"0110111111",
		"0110111001",
		"0110110100",
		"0110101111",
		"0110101010",
		"0110100101",
		"0110100000",
		"0110011011",
		"0110010110",
		"0110010010",
		"0110001101",
		"0110001000",
		"0110000100",
		"0110000000",
		"0101111011",
		"0101110111",
		"0101110011",
		"0101101111",
		"0101101011",
		"0101100111",
		"0101100011",
		"0101011111",
		"0101011011",
		"0101011000",
		"0101010100",
		"0101010001",
		"0101001101",
		"0101001010",
		"0101000110",
		"0101000011",
		"0100111111",
		"0100111100",
		"0100111001",
		"0100110110",
		"0100110011",
		"0100110000",
		"0100101101",
		"0100101010",
		"0100100111",
		"0100100100",
		"0100100001",
		"0100011110",
		"0100011011",
		"0100011001",
		"0100010110",
		"0100010011",
		"0100010001",
		"0100001110",
		"0100001100",
		"0100001001",
		"0100000111",
		"0100000100",
		"0100000010",
		"0011111111",
		"0011111101",
		"0011111011",
		"0011111000",
		"0011110110",
		"0011110100",
		"0011110010",
		"0011110000",
		"0011101101",
		"0011101011",
		"0011101001",
		"0011100111",
		"0011100101",
		"0011100011",
		"0011100001",
		"0011011111",
		"0011011101",
		"0011011100",
		"0011011010",
		"0011011000",
		"0011010110",
		"0011010100",
		"0011010010",
		"0011010001",
		"0011001111",
		"0011001101",
		"0011001100",
		"0011001010",
		"0011001000",
		"0011000111",
		"0011000101",
		"0011000011",
		"0011000010",
		"0011000000",
		"0010111111",
		"0010111101",
		"0010111100",
		"0010111010",
		"0010111001"
	);
begin
	data <= "1"&rom(to_integer(unsigned(addr)))&"000";
end architecture;