library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity LUT_C0_reci_sqrt_1_2 is
	generic(
		word_bits	:natural:=25;
		bus_bits	:natural:=29;
		add_bits	:natural:=7
	);
	port(
		addr		:in std_logic_vector(add_bits-1 downto 0);
		data		:out std_logic_vector(bus_bits-1 downto 0)
	);
end entity;

architecture behav of LUT_C0_reci_sqrt_1_2 is
	type storage is array (0 to 2**add_bits-1) of std_logic_vector(word_bits-1 downto 0);
	signal rom:storage:=(
		"1111111111111111111111111",
		"1111111000000010111110101",
		"1111110000001011110110000",
		"1111101000011010011110111",
		"1111100000101110110010000",
		"1111011001001000101000111",
		"1111010001100111111100100",
		"1111001010001100100110110",
		"1111000010110110100001000",
		"1110111011100101100101011",
		"1110110100011001101101110",
		"1110101101010010110100010",
		"1110100110010000110011011",
		"1110011111010011100101010",
		"1110011000011011000100110",
		"1110010001100111001100100",
		"1110001010110111110111011",
		"1110000100001101000000010",
		"1101111101100110100010011",
		"1101110111000100011000110",
		"1101110000100110011110111",
		"1101101010001100110000001",
		"1101100011110111001000000",
		"1101011101100101100010010",
		"1101010111010111111010100",
		"1101010001001110001100110",
		"1101001011001000010100110",
		"1101000101000110001110101",
		"1100111111000111110110100",
		"1100111001001101001000100",
		"1100110011010110000001000",
		"1100101101100010011100011",
		"1100100111110010010111000",
		"1100100010000101101101100",
		"1100011100011100011100011",
		"1100010110110110100000011",
		"1100010001010011110110001",
		"1100001011110100011010101",
		"1100000110011000001010110",
		"1100000000111111000011010",
		"1011111011101001000001010",
		"1011110110010110000001111",
		"1011110001000110000010010",
		"1011101011111000111111100",
		"1011100110101110110110111",
		"1011100001100111100101101",
		"1011011100100011001001011",
		"1011010111100001011111010",
		"1011010010100010100100111",
		"1011001101100110010111101",
		"1011001000101100110101010",
		"1011000011110101111011010",
		"1010111111000001100111010",
		"1010111010001111110111001",
		"1010110101100000101000011",
		"1010110000110011111001000",
		"1010101100001001100110101",
		"1010100111100001101111011",
		"1010100010111100010001000",
		"1010011110011001001001011",
		"1010011001111000010110110",
		"1010010101011001110111000",
		"1010010000111101101000001",
		"1010001100100011101000010",
		"1010001000001011110101101",
		"1010000011110110001110011",
		"1001111111100010110000110",
		"1001111011010001011010110",
		"1001110111000010001010111",
		"1001110010110100111111011",
		"1001101110101001110110100",
		"1001101010100000101110110",
		"1001100110011001100110011",
		"1001100010010100011011110",
		"1001011110010001001101100",
		"1001011010001111111001111",
		"1001010110010000011111101",
		"1001010010010010111101000",
		"1001001110010111010000110",
		"1001001010011101011001011",
		"1001000110100101010101100",
		"1001000010101111000011101",
		"1000111110111010100010100",
		"1000111011000111110000110",
		"1000110111010110101101000",
		"1000110011100111010110001",
		"1000101111111001101010101",
		"1000101100001101101001100",
		"1000101000100011010001011",
		"1000100100111010100001000",
		"1000100001010011010111011",
		"1000011101101101110011000",
		"1000011010001001110011000",
		"1000010110100111010110010",
		"1000010011000110011011011",
		"1000001111100111000001100",
		"1000001100001001000111100",
		"1000001000101100101100010",
		"1000000101010001101110111",
		"1000000001111000001110000",
		"0111111110100000001000111",
		"0111111011001001011110100",
		"0111110111110100001101110",
		"0111110100100000010101110",
		"0111110001001101110101100",
		"0111101101111100101100001",
		"0111101010101100111000101",
		"0111100111011110011010001",
		"0111100100010001001111101",
		"0111100001000101011000011",
		"0111011101111010110011011",
		"0111011010110001011111111",
		"0111010111101001011101000",
		"0111010100100010101001111",
		"0111010001011101000101110",
		"0111001110011000101111110",
		"0111001011010101100111000",
		"0111001000010011101010111",
		"0111000101010010111010011",
		"0111000010010011010101000",
		"0110111111010100111001111",
		"0110111100010111101000001",
		"0110111001011011011111010",
		"0110110110100000011110010",
		"0110110011100110100100110",
		"0110110000101101110001110",
		"0110101101110110000100101",
		"0110101010111111011100111"
	);
begin
	data <= "001"&rom(to_integer(unsigned(addr)))&"0";
end architecture;