library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity LUT_C1_reci_sqrt_2_4 is
	generic(
		word_bits	:natural:=15;
		bus_bits	:natural:=20;
		add_bits	:natural:=7
	);
	port(
		addr		:in std_logic_vector(add_bits-1 downto 0);
		data		:out std_logic_vector(bus_bits-1 downto 0)
	);
end entity;

architecture behav of LUT_C1_reci_sqrt_2_4 is
	type storage is array (0 to 2**add_bits-1) of std_logic_vector(word_bits-1 downto 0);
	signal rom:storage:=(
		"101101010000001",
		"101100101110101",
		"101100001101101",
		"101011101101010",
		"101011001101100",
		"101010101110011",
		"101010001111111",
		"101001110001111",
		"101001010100011",
		"101000110111100",
		"101000011011001",
		"100111111111010",
		"100111100011111",
		"100111001001000",
		"100110101110101",
		"100110010100101",
		"100101111011001",
		"100101100010001",
		"100101001001100",
		"100100110001010",
		"100100011001011",
		"100100000010000",
		"100011101011000",
		"100011010100011",
		"100010111110001",
		"100010101000001",
		"100010010010101",
		"100001111101011",
		"100001101000100",
		"100001010100000",
		"100000111111111",
		"100000101011111",
		"100000011000011",
		"100000000101000",
		"011111110010001",
		"011111011111011",
		"011111001101000",
		"011110111010111",
		"011110101001000",
		"011110010111011",
		"011110000110001",
		"011101110101000",
		"011101100100010",
		"011101010011101",
		"011101000011010",
		"011100110011010",
		"011100100011011",
		"011100010011101",
		"011100000100010",
		"011011110101001",
		"011011100110001",
		"011011010111010",
		"011011001000110",
		"011010111010011",
		"011010101100001",
		"011010011110010",
		"011010010000011",
		"011010000010110",
		"011001110101011",
		"011001101000001",
		"011001011011000",
		"011001001110001",
		"011001000001011",
		"011000110100111",
		"011000101000100",
		"011000011100010",
		"011000010000001",
		"011000000100010",
		"010111111000100",
		"010111101100111",
		"010111100001011",
		"010111010110000",
		"010111001010111",
		"010110111111110",
		"010110110100111",
		"010110101010001",
		"010110011111011",
		"010110010100111",
		"010110001010100",
		"010110000000010",
		"010101110110001",
		"010101101100001",
		"010101100010001",
		"010101011000011",
		"010101001110110",
		"010101000101001",
		"010100111011110",
		"010100110010011",
		"010100101001001",
		"010100100000000",
		"010100010111000",
		"010100001110001",
		"010100000101010",
		"010011111100101",
		"010011110100000",
		"010011101011100",
		"010011100011000",
		"010011011010101",
		"010011010010100",
		"010011001010010",
		"010011000010010",
		"010010111010010",
		"010010110010011",
		"010010101010101",
		"010010100010111",
		"010010011011010",
		"010010010011101",
		"010010001100010",
		"010010000100111",
		"010001111101100",
		"010001110110010",
		"010001101111001",
		"010001101000000",
		"010001100001000",
		"010001011010001",
		"010001010011010",
		"010001001100011",
		"010001000101101",
		"010000111111000",
		"010000111000011",
		"010000110001111",
		"010000101011011",
		"010000100101000",
		"010000011110101",
		"010000011000011",
		"010000010010010",
		"010000001100000",
		"010000000110000"
	);
begin
	data <= "100"&rom(to_integer(unsigned(addr)))&"00";
end architecture;