library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity LUT_C0_reci is
	generic(
		word_bits	:natural:=25;
		bus_bits	:natural:=29;
		add_bits	:natural:=7
	);
	port(
		addr		:in std_logic_vector(add_bits-1 downto 0);
		data		:out std_logic_vector(bus_bits-1 downto 0)
	);
end entity;

architecture behav of LUT_C0_reci is
	type storage is array (0 to 2**add_bits-1) of std_logic_vector(word_bits-1 downto 0);
	signal rom:storage:=(
		"1111111111111111111111111",
		"1111110000000111111011111",
		"1111100000011111100000011",
		"1111010001000110010110010",
		"1111000001111100000111101",
		"1110110011000000011110101",
		"1110100100010011000110100",
		"1110010101110011101011000",
		"1110000111100001111000010",
		"1101111001011101011011011",
		"1101101011100110000001110",
		"1101011101111011011001001",
		"1101010000011101010000010",
		"1101000011001011010110001",
		"1100110110000101011010000",
		"1100101001001011001100000",
		"1100011100011100011100010",
		"1100001111111000111011111",
		"1100000011100000011011111",
		"1011110111010010101110000",
		"1011101011001111100100010",
		"1011011111010110110000111",
		"1011010011101000000110110",
		"1011001000000011011000111",
		"1010111100101000011010111",
		"1010110001010111000000010",
		"1010100110001110111101011",
		"1010011011010000000110100",
		"1010010000011010010000010",
		"1010000101101101001111110",
		"1001111011001000111010010",
		"1001110000101101000101001",
		"1001100110011001100110010",
		"1001011100001110010011110",
		"1001010010001011000011111",
		"1001001000001111101101000",
		"1000111110011100000110001",
		"1000110100110000000110001",
		"1000101011001011100100001",
		"1000100001101110010111101",
		"1000011000011000011000010",
		"1000001111001001011101111",
		"1000000110000001100000010",
		"0111111101000000010111111",
		"0111110100000101111100111",
		"0111101011010010001000000",
		"0111100010100100110001111",
		"0111011001111101110011100",
		"0111010001011101000101110",
		"0111001001000010100001111",
		"0111000000101110000001011",
		"0110111000011111011101101",
		"0110110000010110110000010",
		"0110101000010011110011001",
		"0110100000010110100000010",
		"0110011000011110110001101",
		"0110010000101100100001010",
		"0110001000111111101001110",
		"0110000001011000000101011",
		"0101111001110101101110110",
		"0101110010011000100000101",
		"0101101011000000010101101",
		"0101100011101101001000101",
		"0101011100011110110100111",
		"0101010101010101010101010",
		"0101001110010000100101000",
		"0101000111010000011111101",
		"0101000000010101000000010",
		"0100111001011110000010100",
		"0100110010101011100010000",
		"0100101011111101011010011",
		"0100100101010011100111100",
		"0100011110101110000101000",
		"0100011000001100101111000",
		"0100010001101111100001100",
		"0100001011010110011000100",
		"0100000101000001010000010",
		"0011111110110000000100111",
		"0011111000100010110010111",
		"0011110010011001010110100",
		"0011101100010011101100010",
		"0011100110010001110000101",
		"0011100000010011100000010",
		"0011011010011000110111110",
		"0011010100100001110011111",
		"0011001110101110010001011",
		"0011001000111110001101001",
		"0011000011010001100100000",
		"0010111101101000010010111",
		"0010111000000010010110111",
		"0010110010011111101101001",
		"0010101101000000010010101",
		"0010100111100100000100101",
		"0010100010001011000000010",
		"0010011100110101000010110",
		"0010010111100010001001101",
		"0010010010010010010010010",
		"0010001101000101011001110",
		"0010000111111011011110000",
		"0010000010110100011100001",
		"0001111101110000010001111",
		"0001111000101110111100111",
		"0001110011110000011010101",
		"0001101110110100101000111",
		"0001101001111011100101100",
		"0001100101000101001101111",
		"0001100000010001100000010",
		"0001011011100000011010001",
		"0001010110110001111001011",
		"0001010010000101111100001",
		"0001001101011100100000010",
		"0001001000110101100011100",
		"0001000100010001000100010",
		"0000111111101111000000010",
		"0000111011001111010101101",
		"0000110110110010000010101",
		"0000110010010111000101001",
		"0000101101111110011011101",
		"0000101001101000000100001",
		"0000100101010011111100111",
		"0000100001000010000100000",
		"0000011100110010011000001",
		"0000011000100100110111010",
		"0000010100011001011111110",
		"0000010000010000010000001",
		"0000001100001001000110110",
		"0000001000000100000010000",
		"0000000100000001000000001"
	);
begin
	data <= "001"&rom(to_integer(unsigned(addr)))&"0";
end architecture;