library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity LUT_C1_exp is
	generic(
		word_bits	:natural:=19;
		bus_bits	:natural:=20;
		add_bits	:natural:=6
	);
	port(
		addr		:in std_logic_vector(add_bits-1 downto 0);
		data		:out std_logic_vector(bus_bits-1 downto 0)
	);
end entity;

architecture behav of LUT_C1_exp is
	type storage is array (0 to 2**add_bits-1) of std_logic_vector(word_bits-1 downto 0);
	signal rom:storage:=(
		"0101100010111000000",
		"0101100110110000000",
		"0101101010101010000",
		"0101101110100110000",
		"0101110010100110000",
		"0101110110101000000",
		"0101111010101101000",
		"0101111110110101000",
		"0110000011000000000",
		"0110000111001110000",
		"0110001011011110000",
		"0110001111110010000",
		"0110010100001001000",
		"0110011000100010000",
		"0110011100111111000",
		"0110100001011111000",
		"0110100110000010000",
		"0110101010101000000",
		"0110101111010001000",
		"0110110011111110000",
		"0110111000101110000",
		"0110111101100001000",
		"0111000010010111000",
		"0111000111010001000",
		"0111001100001110000",
		"0111010001001111000",
		"0111010110010011000",
		"0111011011011011000",
		"0111100000100110000",
		"0111100101110101000",
		"0111101011001000000",
		"0111110000011110000",
		"0111110101111000000",
		"0111111011010110000",
		"1000000000111000000",
		"1000000110011101000",
		"1000001100000110000",
		"1000010001110100000",
		"1000010111100101000",
		"1000011101011010000",
		"1000100011010011000",
		"1000101001010001000",
		"1000101111010010000",
		"1000110101011000000",
		"1000111011100010000",
		"1001000001110001000",
		"1001001000000011000",
		"1001001110011010000",
		"1001010100110110000",
		"1001011011010110000",
		"1001100001111010000",
		"1001101000100011000",
		"1001101111010001000",
		"1001110110000011000",
		"1001111100111010000",
		"1010000011110110000",
		"1010001010110111000",
		"1010010001111101000",
		"1010011001000111000",
		"1010100000010111000",
		"1010100111101011000",
		"1010101111000101000",
		"1010110110100100000",
		"1010111110001000000"
	);
begin
	data <= "0"&rom(to_integer(unsigned(addr)));
end architecture;