library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity LUT_C1_ln2e0 is
	generic(
		word_bits	:natural:=18;
		bus_bits	:natural:=20;
		add_bits	:natural:=6
	);
	port(
		addr		:in std_logic_vector(add_bits-1 downto 0);
		data		:out std_logic_vector(bus_bits-1 downto 0)
	);
end entity;

architecture behav of LUT_C1_ln2e0 is
	type storage is array (0 to 2**add_bits-1) of std_logic_vector(word_bits-1 downto 0);
	signal rom:storage:=(
		"101110001010011000",
		"101101001101111000",
		"101100010011100000",
		"101011011011000000",
		"101010100100011000",
		"101001101111101000",
		"101000111100100000",
		"101000001011000000",
		"100111011011001000",
		"100110101100101000",
		"100101111111101000",
		"100101010011111000",
		"100100101001100000",
		"100100000000011000",
		"100011011000100000",
		"100010110001110000",
		"100010001100000000",
		"100001100111011000",
		"100001000011110000",
		"100000100001001000",
		"011111111111100000",
		"011111011110101000",
		"011110111110110000",
		"011110011111101000",
		"011110000001011000",
		"011101100011111000",
		"011101000111001000",
		"011100101011001000",
		"011100001111110000",
		"011011110101000000",
		"011011011011000000",
		"011011000001101000",
		"011010101000111000",
		"011010010000101000",
		"011001111001000000",
		"011001100010000000",
		"011001001011011000",
		"011000110101011000",
		"011000011111111000",
		"011000001010110000",
		"010111110110001000",
		"010111100010000000",
		"010111001110011000",
		"010110111011000000",
		"010110101000001000",
		"010110010101110000",
		"010110000011101000",
		"010101110001111000",
		"010101100000101000",
		"010101001111101000",
		"010100111111000000",
		"010100101110101000",
		"010100011110101000",
		"010100001111000000",
		"010011111111101000",
		"010011110000101000",
		"010011100001111000",
		"010011010011011000",
		"010011000101001000",
		"010010110111010000",
		"010010101001100000",
		"010010011100001000",
		"010010001110111000",
		"010010000010000000"
	);
begin
	data <= "10"&rom(to_integer(unsigned(addr)));
end architecture;