library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity LUT_C2_reci_sqrt_1_2 is
	generic(
		word_bits	:natural:=12;
		bus_bits	:natural:=14;
		add_bits	:natural:=7
	);
	port(
		addr		:in std_logic_vector(add_bits-1 downto 0);
		data		:out std_logic_vector(bus_bits-1 downto 0)
	);
end entity;

architecture behav of LUT_C2_reci_sqrt_1_2 is
	type storage is array (0 to 2**add_bits-1) of std_logic_vector(word_bits-1 downto 0);
	signal rom:storage:=(
		"101111100000",
		"101110100000",
		"101101101000",
		"101100110000",
		"101100000000",
		"101011001000",
		"101010011000",
		"101001101000",
		"101000110000",
		"101000001000",
		"100111011000",
		"100110101000",
		"100110000000",
		"100101010000",
		"100100101000",
		"100100000000",
		"100011011000",
		"100010110000",
		"100010010000",
		"100001101000",
		"100001000000",
		"100000100000",
		"100000000000",
		"011111011000",
		"011110111000",
		"011110011000",
		"011101111000",
		"011101100000",
		"011101000000",
		"011100100000",
		"011100001000",
		"011011101000",
		"011011010000",
		"011010110000",
		"011010011000",
		"011010000000",
		"011001101000",
		"011001010000",
		"011000110000",
		"011000100000",
		"011000001000",
		"010111110000",
		"010111011000",
		"010111000000",
		"010110110000",
		"010110011000",
		"010110000000",
		"010101110000",
		"010101011000",
		"010101001000",
		"010100111000",
		"010100100000",
		"010100010000",
		"010100000000",
		"010011110000",
		"010011100000",
		"010011001000",
		"010010111000",
		"010010101000",
		"010010011000",
		"010010001000",
		"010001111000",
		"010001110000",
		"010001100000",
		"010001010000",
		"010001000000",
		"010000110000",
		"010000101000",
		"010000011000",
		"010000001000",
		"010000000000",
		"001111110000",
		"001111101000",
		"001111011000",
		"001111001000",
		"001111000000",
		"001110111000",
		"001110101000",
		"001110100000",
		"001110010000",
		"001110001000",
		"001110000000",
		"001101110000",
		"001101101000",
		"001101100000",
		"001101010000",
		"001101001000",
		"001101000000",
		"001100111000",
		"001100110000",
		"001100100000",
		"001100011000",
		"001100010000",
		"001100001000",
		"001100000000",
		"001011111000",
		"001011110000",
		"001011101000",
		"001011100000",
		"001011011000",
		"001011010000",
		"001011001000",
		"001011000000",
		"001010111000",
		"001010110000",
		"001010101000",
		"001010100000",
		"001010011000",
		"001010010000",
		"001010001000",
		"001010001000",
		"001010000000",
		"001001111000",
		"001001110000",
		"001001101000",
		"001001100000",
		"001001100000",
		"001001011000",
		"001001010000",
		"001001001000",
		"001001001000",
		"001001000000",
		"001000111000",
		"001000110000",
		"001000110000",
		"001000101000",
		"001000100000",
		"001000100000"
	);
begin
	data <= "00"&rom(to_integer(unsigned(addr)));
end architecture;