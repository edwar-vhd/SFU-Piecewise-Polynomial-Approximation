library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity LUT_C1_sin is
	generic(
		word_bits	:natural:=19;
		bus_bits	:natural:=20;
		add_bits	:natural:=6
	);
	port(
		addr		:in std_logic_vector(add_bits-1 downto 0);
		data		:out std_logic_vector(bus_bits-1 downto 0)
	);
end entity;

architecture behav of LUT_C1_sin is
	type storage is array (0 to 2**add_bits-1) of std_logic_vector(word_bits-1 downto 0);
	signal rom:storage:=(
		"1000000000000000101",
		"0111111111111100101",
		"0111111111110000110",
		"0111111111011100110",
		"0111111111000000110",
		"0111111110011100110",
		"0111111101110000110",
		"0111111100111100111",
		"0111111100000001000",
		"0111111010111101010",
		"0111111001110001100",
		"0111111000011101111",
		"0111110111000010011",
		"0111110101011111000",
		"0111110011110011110",
		"0111110010000000110",
		"0111110000000110000",
		"0111101110000011100",
		"0111101011111001001",
		"0111101001100111010",
		"0111100111001101101",
		"0111100100101100011",
		"0111100010000011101",
		"0111011111010011011",
		"0111011100011011100",
		"0111011001011100010",
		"0111010110010101101",
		"0111010011000111101",
		"0111001111110010011",
		"0111001100010101110",
		"0111001000110010000",
		"0111000101000111001",
		"0111000001010101010",
		"0110111101011100010",
		"0110111001011100011",
		"0110110101010101100",
		"0110110001000111111",
		"0110101100110011011",
		"0110101000011000010",
		"0110100011110110100",
		"0110011111001110001",
		"0110011010011111011",
		"0110010101101010001",
		"0110010000101110101",
		"0110001011101100110",
		"0110000110100100110",
		"0110000001010110101",
		"0101111100000010100",
		"0101110110101000100",
		"0101110001001000100",
		"0101101011100010111",
		"0101100101110111100",
		"0101100000000110100",
		"0101011010010000001",
		"0101010100010100010",
		"0101001110010011000",
		"0101001000001100101",
		"0101000010000001000",
		"0100111011110000100",
		"0100110101011011000",
		"0100101111000000101",
		"0100101000100001101",
		"0100100001111101111",
		"0100011011010101101"
	);
begin
	data <= "0"&rom(to_integer(unsigned(addr)));
end architecture;