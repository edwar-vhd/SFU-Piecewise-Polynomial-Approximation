library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity LUT_C1_reci_sqrt_1_2 is
	generic(
		word_bits	:natural:=15;
		bus_bits	:natural:=20;
		add_bits	:natural:=7
	);
	port(
		addr		:in std_logic_vector(add_bits-1 downto 0);
		data		:out std_logic_vector(bus_bits-1 downto 0)
	);
end entity;

architecture behav of LUT_C1_reci_sqrt_1_2 is
	type storage is array (0 to 2**add_bits-1) of std_logic_vector(word_bits-1 downto 0);
	signal rom:storage:=(
		"111111111111111",
		"111111010000011",
		"111110100001110",
		"111101110100000",
		"111101000111001",
		"111100011011001",
		"111011101111111",
		"111011000101100",
		"111010011011111",
		"111001110011000",
		"111001001010111",
		"111000100011011",
		"110111111100110",
		"110111010110101",
		"110110110001011",
		"110110001100101",
		"110101101000100",
		"110101000101001",
		"110100100010010",
		"110100000000000",
		"110011011110011",
		"110010111101010",
		"110010011100101",
		"110001111100101",
		"110001011101001",
		"110000111110001",
		"110000011111110",
		"110000000001110",
		"101111100100010",
		"101111000111001",
		"101110101010101",
		"101110001110100",
		"101101110010110",
		"101101010111100",
		"101100111100101",
		"101100100010010",
		"101100001000010",
		"101011101110100",
		"101011010101010",
		"101010111100011",
		"101010100011111",
		"101010001011110",
		"101001110100000",
		"101001011100100",
		"101001000101100",
		"101000101110110",
		"101000011000010",
		"101000000010001",
		"100111101100011",
		"100111010110111",
		"100111000001101",
		"100110101100110",
		"100110011000001",
		"100110000011110",
		"100101101111110",
		"100101011100000",
		"100101001000100",
		"100100110101010",
		"100100100010010",
		"100100001111100",
		"100011111101000",
		"100011101010110",
		"100011011000110",
		"100011000111000",
		"100010110101100",
		"100010100100010",
		"100010010011001",
		"100010000010010",
		"100001110001101",
		"100001100001001",
		"100001010000111",
		"100001000000111",
		"100000110001001",
		"100000100001100",
		"100000010010000",
		"100000000010110",
		"011111110011110",
		"011111100100111",
		"011111010110001",
		"011111000111101",
		"011110111001010",
		"011110101011001",
		"011110011101001",
		"011110001111010",
		"011110000001100",
		"011101110100000",
		"011101100110101",
		"011101011001100",
		"011101001100011",
		"011100111111100",
		"011100110010110",
		"011100100110001",
		"011100011001110",
		"011100001101011",
		"011100000001010",
		"011011110101001",
		"011011101001010",
		"011011011101100",
		"011011010001110",
		"011011000110010",
		"011010111010111",
		"011010101111101",
		"011010100100100",
		"011010011001011",
		"011010001110100",
		"011010000011110",
		"011001111001000",
		"011001101110100",
		"011001100100000",
		"011001011001101",
		"011001001111011",
		"011001000101010",
		"011000111011010",
		"011000110001011",
		"011000100111100",
		"011000011101111",
		"011000010100010",
		"011000001010110",
		"011000000001010",
		"010111111000000",
		"010111101110110",
		"010111100101101",
		"010111011100100",
		"010111010011101",
		"010111001010110",
		"010111000001111",
		"010110111001010",
		"010110110000101"
	);
begin
	data <= "100"&rom(to_integer(unsigned(addr)))&"00";
end architecture;