library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity LUT_C0_reci_sqrt_2_4 is
	generic(
		word_bits	:natural:=25;
		bus_bits	:natural:=29;
		add_bits	:natural:=7
	);
	port(
		addr		:in std_logic_vector(add_bits-1 downto 0);
		data		:out std_logic_vector(bus_bits-1 downto 0)
	);
end entity;

architecture behav of LUT_C0_reci_sqrt_2_4 is
	type storage is array (0 to 2**add_bits-1) of std_logic_vector(word_bits-1 downto 0);
	signal rom:storage:=(
		"1101010000010011110011000",
		"1101000101000011111011110",
		"1100111001111100011001010",
		"1100101110111101000001010",
		"1100100100000101101001100",
		"1100011001010110001000110",
		"1100001110101110010101100",
		"1100000100001110000110100",
		"1011111001110101010011000",
		"1011101111100011110010010",
		"1011100101011001011011100",
		"1011011011010110000111000",
		"1011010001011001101100010",
		"1011000111100100000011100",
		"1010111101110101000101010",
		"1010110100001100101010000",
		"1010101010101010101010100",
		"1010100001001110111111100",
		"1010010111111001100010000",
		"1010001110101010001011100",
		"1010000101100000110101000",
		"1001111100011101011000100",
		"1001110011011111101111100",
		"1001101010100111110011110",
		"1001100001110101011111010",
		"1001011001001000101100000",
		"1001010000100001010100100",
		"1001000111111111010011010",
		"1000111111100010100010010",
		"1000110111001010111100110",
		"1000101110111000011101000",
		"1000100110101010111110000",
		"1000011110100010011011000",
		"1000010110011110101110110",
		"1000001110011111110100100",
		"1000000110100101100111110",
		"0111111110110000000011100",
		"0111110110111111000011110",
		"0111101111010010100011110",
		"0111100111101010011111100",
		"0111100000000110110010100",
		"0111011000100111011000100",
		"0111010001001100001101110",
		"0111001001110101001110000",
		"0111000010100010010101110",
		"0110111011010011100000110",
		"0110110100001000101011100",
		"0110101101000001110010100",
		"0110100101111110110001110",
		"0110011110111111100110000",
		"0110011000000100001100000",
		"0110010001001100011111110",
		"0110001010011000011110110",
		"0110000011101000000101000",
		"0101111100111011001111110",
		"0101110110010001111011110",
		"0101101111101100000110000",
		"0101101001001001101011100",
		"0101100010101010101001010",
		"0101011100001110111100010",
		"0101010101110110100001110",
		"0101001111100001010111000",
		"0101001001001111011001010",
		"0101000011000000100101110",
		"0100111100110100111010000",
		"0100110110101100010011010",
		"0100110000100110101111010",
		"0100101010100100001011000",
		"0100100100100100100100100",
		"0100011110100111111001000",
		"0100011000101110000110100",
		"0100010010110111001010010",
		"0100001101000011000010100",
		"0100000111010001101100100",
		"0100000001100011000110010",
		"0011111011110111001101100",
		"0011110110001110000000100",
		"0011110000100111011100100",
		"0011101011000011100000000",
		"0011100101100010001000110",
		"0011100000000011010100110",
		"0011011010100111000010010",
		"0011010101001101001111000",
		"0011001111110101111001010",
		"0011001010100000111111010",
		"0011000101001110011111000",
		"0010111111111110010110110",
		"0010111010110000100101000",
		"0010110101100101000111100",
		"0010110000011011111101000",
		"0010101011010101000011100",
		"0010100110010000011001100",
		"0010100001001101111101010",
		"0010011100001101101101010",
		"0010010111001111101000000",
		"0010010010010011101011110",
		"0010001101011001110111000",
		"0010001000100010001000100",
		"0010000011101100011110010",
		"0001111110111000110111010",
		"0001111010000111010010000",
		"0001110101010111101101000",
		"0001110000101010000110110",
		"0001101011111110011110000",
		"0001100111010100110001100",
		"0001100010101100111111100",
		"0001011110000111000111010",
		"0001011001100011000111000",
		"0001010101000000111101110",
		"0001010000100000101010010",
		"0001001100000010001011000",
		"0001000111100101011111000",
		"0001000011001010100101000",
		"0000111110110001011011110",
		"0000111010011010000010010",
		"0000110110000100010111010",
		"0000110001110000011001100",
		"0000101101011110001000000",
		"0000101001001101100001110",
		"0000100100111110100101100",
		"0000100000110001010010000",
		"0000011100100101100110110",
		"0000011000011011100010010",
		"0000010100010011000011110",
		"0000010000001100001010000",
		"0000001100000110110100010",
		"0000001000000011000001010",
		"0000000100000000110000000"
	);
begin
	data <= "0010"&rom(to_integer(unsigned(addr)));
end architecture;