library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity LUT_C2_sqrt_2_4 is
	generic(
		word_bits	:natural:=11;
		bus_bits	:natural:=14;
		add_bits	:natural:=6
	);
	port(
		addr		:in std_logic_vector(add_bits-1 downto 0);
		data		:out std_logic_vector(bus_bits-1 downto 0)
	);
end entity;

architecture behav of LUT_C2_sqrt_2_4 is
	type storage is array (0 to 2**add_bits-1) of std_logic_vector(word_bits-1 downto 0);
	signal rom:storage:=(
		"10110010100",
		"10101110100",
		"10101010100",
		"10100111000",
		"10100011000",
		"10011111100",
		"10011100100",
		"10011001000",
		"10010110000",
		"10010011000",
		"10010000000",
		"10001101000",
		"10001010100",
		"10000111100",
		"10000101000",
		"10000010100",
		"10000000000",
		"01111101100",
		"01111011100",
		"01111001000",
		"01110111000",
		"01110101000",
		"01110011000",
		"01110001000",
		"01101111000",
		"01101101000",
		"01101011100",
		"01101001100",
		"01101000000",
		"01100110100",
		"01100100100",
		"01100011000",
		"01100001100",
		"01100000000",
		"01011110100",
		"01011101000",
		"01011011100",
		"01011010100",
		"01011001000",
		"01011000000",
		"01010110100",
		"01010101100",
		"01010100000",
		"01010011000",
		"01010010000",
		"01010000100",
		"01001111100",
		"01001110100",
		"01001101100",
		"01001100100",
		"01001011100",
		"01001010100",
		"01001001100",
		"01001000100",
		"01000111100",
		"01000110100",
		"01000110000",
		"01000101000",
		"01000100000",
		"01000011100",
		"01000010100",
		"01000001100",
		"01000001000",
		"01000000000"
	);
begin
	data <= "100"&rom(to_integer(unsigned(addr)));
end architecture;